magic
tech sky130A
magscale 1 2
timestamp 1731174374
<< metal4 >>
rect -10294 4039 -7196 4080
rect -10294 1561 -7452 4039
rect -7216 1561 -7196 4039
rect -10294 1520 -7196 1561
rect -6796 4039 -3698 4080
rect -6796 1561 -3954 4039
rect -3718 1561 -3698 4039
rect -6796 1520 -3698 1561
rect -3298 4039 -200 4080
rect -3298 1561 -456 4039
rect -220 1561 -200 4039
rect -3298 1520 -200 1561
rect 200 4039 3298 4080
rect 200 1561 3042 4039
rect 3278 1561 3298 4039
rect 200 1520 3298 1561
rect 3698 4039 6796 4080
rect 3698 1561 6540 4039
rect 6776 1561 6796 4039
rect 3698 1520 6796 1561
rect 7196 4039 10294 4080
rect 7196 1561 10038 4039
rect 10274 1561 10294 4039
rect 7196 1520 10294 1561
rect -10294 1239 -7196 1280
rect -10294 -1239 -7452 1239
rect -7216 -1239 -7196 1239
rect -10294 -1280 -7196 -1239
rect -6796 1239 -3698 1280
rect -6796 -1239 -3954 1239
rect -3718 -1239 -3698 1239
rect -6796 -1280 -3698 -1239
rect -3298 1239 -200 1280
rect -3298 -1239 -456 1239
rect -220 -1239 -200 1239
rect -3298 -1280 -200 -1239
rect 200 1239 3298 1280
rect 200 -1239 3042 1239
rect 3278 -1239 3298 1239
rect 200 -1280 3298 -1239
rect 3698 1239 6796 1280
rect 3698 -1239 6540 1239
rect 6776 -1239 6796 1239
rect 3698 -1280 6796 -1239
rect 7196 1239 10294 1280
rect 7196 -1239 10038 1239
rect 10274 -1239 10294 1239
rect 7196 -1280 10294 -1239
rect -10294 -1561 -7196 -1520
rect -10294 -4039 -7452 -1561
rect -7216 -4039 -7196 -1561
rect -10294 -4080 -7196 -4039
rect -6796 -1561 -3698 -1520
rect -6796 -4039 -3954 -1561
rect -3718 -4039 -3698 -1561
rect -6796 -4080 -3698 -4039
rect -3298 -1561 -200 -1520
rect -3298 -4039 -456 -1561
rect -220 -4039 -200 -1561
rect -3298 -4080 -200 -4039
rect 200 -1561 3298 -1520
rect 200 -4039 3042 -1561
rect 3278 -4039 3298 -1561
rect 200 -4080 3298 -4039
rect 3698 -1561 6796 -1520
rect 3698 -4039 6540 -1561
rect 6776 -4039 6796 -1561
rect 3698 -4080 6796 -4039
rect 7196 -1561 10294 -1520
rect 7196 -4039 10038 -1561
rect 10274 -4039 10294 -1561
rect 7196 -4080 10294 -4039
<< via4 >>
rect -7452 1561 -7216 4039
rect -3954 1561 -3718 4039
rect -456 1561 -220 4039
rect 3042 1561 3278 4039
rect 6540 1561 6776 4039
rect 10038 1561 10274 4039
rect -7452 -1239 -7216 1239
rect -3954 -1239 -3718 1239
rect -456 -1239 -220 1239
rect 3042 -1239 3278 1239
rect 6540 -1239 6776 1239
rect 10038 -1239 10274 1239
rect -7452 -4039 -7216 -1561
rect -3954 -4039 -3718 -1561
rect -456 -4039 -220 -1561
rect 3042 -4039 3278 -1561
rect 6540 -4039 6776 -1561
rect 10038 -4039 10274 -1561
<< mimcap2 >>
rect -10214 3960 -7814 4000
rect -10214 1640 -10174 3960
rect -7854 1640 -7814 3960
rect -10214 1600 -7814 1640
rect -6716 3960 -4316 4000
rect -6716 1640 -6676 3960
rect -4356 1640 -4316 3960
rect -6716 1600 -4316 1640
rect -3218 3960 -818 4000
rect -3218 1640 -3178 3960
rect -858 1640 -818 3960
rect -3218 1600 -818 1640
rect 280 3960 2680 4000
rect 280 1640 320 3960
rect 2640 1640 2680 3960
rect 280 1600 2680 1640
rect 3778 3960 6178 4000
rect 3778 1640 3818 3960
rect 6138 1640 6178 3960
rect 3778 1600 6178 1640
rect 7276 3960 9676 4000
rect 7276 1640 7316 3960
rect 9636 1640 9676 3960
rect 7276 1600 9676 1640
rect -10214 1160 -7814 1200
rect -10214 -1160 -10174 1160
rect -7854 -1160 -7814 1160
rect -10214 -1200 -7814 -1160
rect -6716 1160 -4316 1200
rect -6716 -1160 -6676 1160
rect -4356 -1160 -4316 1160
rect -6716 -1200 -4316 -1160
rect -3218 1160 -818 1200
rect -3218 -1160 -3178 1160
rect -858 -1160 -818 1160
rect -3218 -1200 -818 -1160
rect 280 1160 2680 1200
rect 280 -1160 320 1160
rect 2640 -1160 2680 1160
rect 280 -1200 2680 -1160
rect 3778 1160 6178 1200
rect 3778 -1160 3818 1160
rect 6138 -1160 6178 1160
rect 3778 -1200 6178 -1160
rect 7276 1160 9676 1200
rect 7276 -1160 7316 1160
rect 9636 -1160 9676 1160
rect 7276 -1200 9676 -1160
rect -10214 -1640 -7814 -1600
rect -10214 -3960 -10174 -1640
rect -7854 -3960 -7814 -1640
rect -10214 -4000 -7814 -3960
rect -6716 -1640 -4316 -1600
rect -6716 -3960 -6676 -1640
rect -4356 -3960 -4316 -1640
rect -6716 -4000 -4316 -3960
rect -3218 -1640 -818 -1600
rect -3218 -3960 -3178 -1640
rect -858 -3960 -818 -1640
rect -3218 -4000 -818 -3960
rect 280 -1640 2680 -1600
rect 280 -3960 320 -1640
rect 2640 -3960 2680 -1640
rect 280 -4000 2680 -3960
rect 3778 -1640 6178 -1600
rect 3778 -3960 3818 -1640
rect 6138 -3960 6178 -1640
rect 3778 -4000 6178 -3960
rect 7276 -1640 9676 -1600
rect 7276 -3960 7316 -1640
rect 9636 -3960 9676 -1640
rect 7276 -4000 9676 -3960
<< mimcap2contact >>
rect -10174 1640 -7854 3960
rect -6676 1640 -4356 3960
rect -3178 1640 -858 3960
rect 320 1640 2640 3960
rect 3818 1640 6138 3960
rect 7316 1640 9636 3960
rect -10174 -1160 -7854 1160
rect -6676 -1160 -4356 1160
rect -3178 -1160 -858 1160
rect 320 -1160 2640 1160
rect 3818 -1160 6138 1160
rect 7316 -1160 9636 1160
rect -10174 -3960 -7854 -1640
rect -6676 -3960 -4356 -1640
rect -3178 -3960 -858 -1640
rect 320 -3960 2640 -1640
rect 3818 -3960 6138 -1640
rect 7316 -3960 9636 -1640
<< metal5 >>
rect -9174 3984 -8854 4200
rect -7494 4039 -7174 4200
rect -10198 3960 -7830 3984
rect -10198 1640 -10174 3960
rect -7854 1640 -7830 3960
rect -10198 1616 -7830 1640
rect -9174 1184 -8854 1616
rect -7494 1561 -7452 4039
rect -7216 1561 -7174 4039
rect -5676 3984 -5356 4200
rect -3996 4039 -3676 4200
rect -6700 3960 -4332 3984
rect -6700 1640 -6676 3960
rect -4356 1640 -4332 3960
rect -6700 1616 -4332 1640
rect -7494 1239 -7174 1561
rect -10198 1160 -7830 1184
rect -10198 -1160 -10174 1160
rect -7854 -1160 -7830 1160
rect -10198 -1184 -7830 -1160
rect -9174 -1616 -8854 -1184
rect -7494 -1239 -7452 1239
rect -7216 -1239 -7174 1239
rect -5676 1184 -5356 1616
rect -3996 1561 -3954 4039
rect -3718 1561 -3676 4039
rect -2178 3984 -1858 4200
rect -498 4039 -178 4200
rect -3202 3960 -834 3984
rect -3202 1640 -3178 3960
rect -858 1640 -834 3960
rect -3202 1616 -834 1640
rect -3996 1239 -3676 1561
rect -6700 1160 -4332 1184
rect -6700 -1160 -6676 1160
rect -4356 -1160 -4332 1160
rect -6700 -1184 -4332 -1160
rect -7494 -1561 -7174 -1239
rect -10198 -1640 -7830 -1616
rect -10198 -3960 -10174 -1640
rect -7854 -3960 -7830 -1640
rect -10198 -3984 -7830 -3960
rect -9174 -4200 -8854 -3984
rect -7494 -4039 -7452 -1561
rect -7216 -4039 -7174 -1561
rect -5676 -1616 -5356 -1184
rect -3996 -1239 -3954 1239
rect -3718 -1239 -3676 1239
rect -2178 1184 -1858 1616
rect -498 1561 -456 4039
rect -220 1561 -178 4039
rect 1320 3984 1640 4200
rect 3000 4039 3320 4200
rect 296 3960 2664 3984
rect 296 1640 320 3960
rect 2640 1640 2664 3960
rect 296 1616 2664 1640
rect -498 1239 -178 1561
rect -3202 1160 -834 1184
rect -3202 -1160 -3178 1160
rect -858 -1160 -834 1160
rect -3202 -1184 -834 -1160
rect -3996 -1561 -3676 -1239
rect -6700 -1640 -4332 -1616
rect -6700 -3960 -6676 -1640
rect -4356 -3960 -4332 -1640
rect -6700 -3984 -4332 -3960
rect -7494 -4200 -7174 -4039
rect -5676 -4200 -5356 -3984
rect -3996 -4039 -3954 -1561
rect -3718 -4039 -3676 -1561
rect -2178 -1616 -1858 -1184
rect -498 -1239 -456 1239
rect -220 -1239 -178 1239
rect 1320 1184 1640 1616
rect 3000 1561 3042 4039
rect 3278 1561 3320 4039
rect 4818 3984 5138 4200
rect 6498 4039 6818 4200
rect 3794 3960 6162 3984
rect 3794 1640 3818 3960
rect 6138 1640 6162 3960
rect 3794 1616 6162 1640
rect 3000 1239 3320 1561
rect 296 1160 2664 1184
rect 296 -1160 320 1160
rect 2640 -1160 2664 1160
rect 296 -1184 2664 -1160
rect -498 -1561 -178 -1239
rect -3202 -1640 -834 -1616
rect -3202 -3960 -3178 -1640
rect -858 -3960 -834 -1640
rect -3202 -3984 -834 -3960
rect -3996 -4200 -3676 -4039
rect -2178 -4200 -1858 -3984
rect -498 -4039 -456 -1561
rect -220 -4039 -178 -1561
rect 1320 -1616 1640 -1184
rect 3000 -1239 3042 1239
rect 3278 -1239 3320 1239
rect 4818 1184 5138 1616
rect 6498 1561 6540 4039
rect 6776 1561 6818 4039
rect 8316 3984 8636 4200
rect 9996 4039 10316 4200
rect 7292 3960 9660 3984
rect 7292 1640 7316 3960
rect 9636 1640 9660 3960
rect 7292 1616 9660 1640
rect 6498 1239 6818 1561
rect 3794 1160 6162 1184
rect 3794 -1160 3818 1160
rect 6138 -1160 6162 1160
rect 3794 -1184 6162 -1160
rect 3000 -1561 3320 -1239
rect 296 -1640 2664 -1616
rect 296 -3960 320 -1640
rect 2640 -3960 2664 -1640
rect 296 -3984 2664 -3960
rect -498 -4200 -178 -4039
rect 1320 -4200 1640 -3984
rect 3000 -4039 3042 -1561
rect 3278 -4039 3320 -1561
rect 4818 -1616 5138 -1184
rect 6498 -1239 6540 1239
rect 6776 -1239 6818 1239
rect 8316 1184 8636 1616
rect 9996 1561 10038 4039
rect 10274 1561 10316 4039
rect 9996 1239 10316 1561
rect 7292 1160 9660 1184
rect 7292 -1160 7316 1160
rect 9636 -1160 9660 1160
rect 7292 -1184 9660 -1160
rect 6498 -1561 6818 -1239
rect 3794 -1640 6162 -1616
rect 3794 -3960 3818 -1640
rect 6138 -3960 6162 -1640
rect 3794 -3984 6162 -3960
rect 3000 -4200 3320 -4039
rect 4818 -4200 5138 -3984
rect 6498 -4039 6540 -1561
rect 6776 -4039 6818 -1561
rect 8316 -1616 8636 -1184
rect 9996 -1239 10038 1239
rect 10274 -1239 10316 1239
rect 9996 -1561 10316 -1239
rect 7292 -1640 9660 -1616
rect 7292 -3960 7316 -1640
rect 9636 -3960 9660 -1640
rect 7292 -3984 9660 -3960
rect 6498 -4200 6818 -4039
rect 8316 -4200 8636 -3984
rect 9996 -4039 10038 -1561
rect 10274 -4039 10316 -1561
rect 9996 -4200 10316 -4039
<< properties >>
string FIXED_BBOX 7196 1520 9756 4080
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 12 l 12 val 297.12 carea 2.00 cperi 0.19 class capacitor nx 6 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
