magic
tech sky130A
magscale 1 2
timestamp 1731176099
<< metal3 >>
rect -8916 4092 -6104 4120
rect -8916 1668 -6188 4092
rect -6124 1668 -6104 4092
rect -8916 1640 -6104 1668
rect -5418 4092 -2606 4120
rect -5418 1668 -2690 4092
rect -2626 1668 -2606 4092
rect -5418 1640 -2606 1668
rect -1920 4092 892 4120
rect -1920 1668 808 4092
rect 872 1668 892 4092
rect -1920 1640 892 1668
rect 1578 4092 4390 4120
rect 1578 1668 4306 4092
rect 4370 1668 4390 4092
rect 1578 1640 4390 1668
rect 5076 4092 7888 4120
rect 5076 1668 7804 4092
rect 7868 1668 7888 4092
rect 5076 1640 7888 1668
rect 8574 4092 11386 4120
rect 8574 1668 11302 4092
rect 11366 1668 11386 4092
rect 8574 1640 11386 1668
rect -8916 1292 -6104 1320
rect -8916 -1132 -6188 1292
rect -6124 -1132 -6104 1292
rect -8916 -1160 -6104 -1132
rect -5418 1292 -2606 1320
rect -5418 -1132 -2690 1292
rect -2626 -1132 -2606 1292
rect -5418 -1160 -2606 -1132
rect -1920 1292 892 1320
rect -1920 -1132 808 1292
rect 872 -1132 892 1292
rect -1920 -1160 892 -1132
rect 1578 1292 4390 1320
rect 1578 -1132 4306 1292
rect 4370 -1132 4390 1292
rect 1578 -1160 4390 -1132
rect 5076 1292 7888 1320
rect 5076 -1132 7804 1292
rect 7868 -1132 7888 1292
rect 5076 -1160 7888 -1132
rect 8574 1292 11386 1320
rect 8574 -1132 11302 1292
rect 11366 -1132 11386 1292
rect 8574 -1160 11386 -1132
rect -8916 -1508 -6104 -1480
rect -8916 -3932 -6188 -1508
rect -6124 -3932 -6104 -1508
rect -8916 -3960 -6104 -3932
rect -5418 -1508 -2606 -1480
rect -5418 -3932 -2690 -1508
rect -2626 -3932 -2606 -1508
rect -5418 -3960 -2606 -3932
rect -1920 -1508 892 -1480
rect -1920 -3932 808 -1508
rect 872 -3932 892 -1508
rect -1920 -3960 892 -3932
rect 1578 -1508 4390 -1480
rect 1578 -3932 4306 -1508
rect 4370 -3932 4390 -1508
rect 1578 -3960 4390 -3932
rect 5076 -1508 7888 -1480
rect 5076 -3932 7804 -1508
rect 7868 -3932 7888 -1508
rect 5076 -3960 7888 -3932
rect 8574 -1508 11386 -1480
rect 8574 -3932 11302 -1508
rect 11366 -3932 11386 -1508
rect 8574 -3960 11386 -3932
<< via3 >>
rect -6188 1668 -6124 4092
rect -2690 1668 -2626 4092
rect 808 1668 872 4092
rect 4306 1668 4370 4092
rect 7804 1668 7868 4092
rect 11302 1668 11366 4092
rect -6188 -1132 -6124 1292
rect -2690 -1132 -2626 1292
rect 808 -1132 872 1292
rect 4306 -1132 4370 1292
rect 7804 -1132 7868 1292
rect 11302 -1132 11366 1292
rect -6188 -3932 -6124 -1508
rect -2690 -3932 -2626 -1508
rect 808 -3932 872 -1508
rect 4306 -3932 4370 -1508
rect 7804 -3932 7868 -1508
rect 11302 -3932 11366 -1508
<< mimcap >>
rect -8876 4040 -6476 4080
rect -8876 1720 -8836 4040
rect -6516 1720 -6476 4040
rect -8876 1680 -6476 1720
rect -5378 4040 -2978 4080
rect -5378 1720 -5338 4040
rect -3018 1720 -2978 4040
rect -5378 1680 -2978 1720
rect -1880 4040 520 4080
rect -1880 1720 -1840 4040
rect 480 1720 520 4040
rect -1880 1680 520 1720
rect 1618 4040 4018 4080
rect 1618 1720 1658 4040
rect 3978 1720 4018 4040
rect 1618 1680 4018 1720
rect 5116 4040 7516 4080
rect 5116 1720 5156 4040
rect 7476 1720 7516 4040
rect 5116 1680 7516 1720
rect 8614 4040 11014 4080
rect 8614 1720 8654 4040
rect 10974 1720 11014 4040
rect 8614 1680 11014 1720
rect -8876 1240 -6476 1280
rect -8876 -1080 -8836 1240
rect -6516 -1080 -6476 1240
rect -8876 -1120 -6476 -1080
rect -5378 1240 -2978 1280
rect -5378 -1080 -5338 1240
rect -3018 -1080 -2978 1240
rect -5378 -1120 -2978 -1080
rect -1880 1240 520 1280
rect -1880 -1080 -1840 1240
rect 480 -1080 520 1240
rect -1880 -1120 520 -1080
rect 1618 1240 4018 1280
rect 1618 -1080 1658 1240
rect 3978 -1080 4018 1240
rect 1618 -1120 4018 -1080
rect 5116 1240 7516 1280
rect 5116 -1080 5156 1240
rect 7476 -1080 7516 1240
rect 5116 -1120 7516 -1080
rect 8614 1240 11014 1280
rect 8614 -1080 8654 1240
rect 10974 -1080 11014 1240
rect 8614 -1120 11014 -1080
rect -8876 -1560 -6476 -1520
rect -8876 -3880 -8836 -1560
rect -6516 -3880 -6476 -1560
rect -8876 -3920 -6476 -3880
rect -5378 -1560 -2978 -1520
rect -5378 -3880 -5338 -1560
rect -3018 -3880 -2978 -1560
rect -5378 -3920 -2978 -3880
rect -1880 -1560 520 -1520
rect -1880 -3880 -1840 -1560
rect 480 -3880 520 -1560
rect -1880 -3920 520 -3880
rect 1618 -1560 4018 -1520
rect 1618 -3880 1658 -1560
rect 3978 -3880 4018 -1560
rect 1618 -3920 4018 -3880
rect 5116 -1560 7516 -1520
rect 5116 -3880 5156 -1560
rect 7476 -3880 7516 -1560
rect 5116 -3920 7516 -3880
rect 8614 -1560 11014 -1520
rect 8614 -3880 8654 -1560
rect 10974 -3880 11014 -1560
rect 8614 -3920 11014 -3880
<< mimcapcontact >>
rect -8836 1720 -6516 4040
rect -5338 1720 -3018 4040
rect -1840 1720 480 4040
rect 1658 1720 3978 4040
rect 5156 1720 7476 4040
rect 8654 1720 10974 4040
rect -8836 -1080 -6516 1240
rect -5338 -1080 -3018 1240
rect -1840 -1080 480 1240
rect 1658 -1080 3978 1240
rect 5156 -1080 7476 1240
rect 8654 -1080 10974 1240
rect -8836 -3880 -6516 -1560
rect -5338 -3880 -3018 -1560
rect -1840 -3880 480 -1560
rect 1658 -3880 3978 -1560
rect 5156 -3880 7476 -1560
rect 8654 -3880 10974 -1560
<< metal4 >>
rect -7728 4041 -7624 4240
rect -6208 4092 -6104 4240
rect -8837 4040 -6515 4041
rect -8837 1720 -8836 4040
rect -6516 1720 -6515 4040
rect -8837 1719 -6515 1720
rect -7728 1241 -7624 1719
rect -6208 1668 -6188 4092
rect -6124 1668 -6104 4092
rect -4230 4041 -4126 4240
rect -2710 4092 -2606 4240
rect -5339 4040 -3017 4041
rect -5339 1720 -5338 4040
rect -3018 1720 -3017 4040
rect -5339 1719 -3017 1720
rect -6208 1292 -6104 1668
rect -8837 1240 -6515 1241
rect -8837 -1080 -8836 1240
rect -6516 -1080 -6515 1240
rect -8837 -1081 -6515 -1080
rect -7728 -1559 -7624 -1081
rect -6208 -1132 -6188 1292
rect -6124 -1132 -6104 1292
rect -4230 1241 -4126 1719
rect -2710 1668 -2690 4092
rect -2626 1668 -2606 4092
rect -732 4041 -628 4240
rect 788 4092 892 4240
rect -1841 4040 481 4041
rect -1841 1720 -1840 4040
rect 480 1720 481 4040
rect -1841 1719 481 1720
rect -2710 1292 -2606 1668
rect -5339 1240 -3017 1241
rect -5339 -1080 -5338 1240
rect -3018 -1080 -3017 1240
rect -5339 -1081 -3017 -1080
rect -6208 -1508 -6104 -1132
rect -8837 -1560 -6515 -1559
rect -8837 -3880 -8836 -1560
rect -6516 -3880 -6515 -1560
rect -8837 -3881 -6515 -3880
rect -7728 -4080 -7624 -3881
rect -6208 -3932 -6188 -1508
rect -6124 -3932 -6104 -1508
rect -4230 -1559 -4126 -1081
rect -2710 -1132 -2690 1292
rect -2626 -1132 -2606 1292
rect -732 1241 -628 1719
rect 788 1668 808 4092
rect 872 1668 892 4092
rect 2766 4041 2870 4240
rect 4286 4092 4390 4240
rect 1657 4040 3979 4041
rect 1657 1720 1658 4040
rect 3978 1720 3979 4040
rect 1657 1719 3979 1720
rect 788 1292 892 1668
rect -1841 1240 481 1241
rect -1841 -1080 -1840 1240
rect 480 -1080 481 1240
rect -1841 -1081 481 -1080
rect -2710 -1508 -2606 -1132
rect -5339 -1560 -3017 -1559
rect -5339 -3880 -5338 -1560
rect -3018 -3880 -3017 -1560
rect -5339 -3881 -3017 -3880
rect -6208 -4080 -6104 -3932
rect -4230 -4080 -4126 -3881
rect -2710 -3932 -2690 -1508
rect -2626 -3932 -2606 -1508
rect -732 -1559 -628 -1081
rect 788 -1132 808 1292
rect 872 -1132 892 1292
rect 2766 1241 2870 1719
rect 4286 1668 4306 4092
rect 4370 1668 4390 4092
rect 6264 4041 6368 4240
rect 7784 4092 7888 4240
rect 5155 4040 7477 4041
rect 5155 1720 5156 4040
rect 7476 1720 7477 4040
rect 5155 1719 7477 1720
rect 4286 1292 4390 1668
rect 1657 1240 3979 1241
rect 1657 -1080 1658 1240
rect 3978 -1080 3979 1240
rect 1657 -1081 3979 -1080
rect 788 -1508 892 -1132
rect -1841 -1560 481 -1559
rect -1841 -3880 -1840 -1560
rect 480 -3880 481 -1560
rect -1841 -3881 481 -3880
rect -2710 -4080 -2606 -3932
rect -732 -4080 -628 -3881
rect 788 -3932 808 -1508
rect 872 -3932 892 -1508
rect 2766 -1559 2870 -1081
rect 4286 -1132 4306 1292
rect 4370 -1132 4390 1292
rect 6264 1241 6368 1719
rect 7784 1668 7804 4092
rect 7868 1668 7888 4092
rect 9762 4041 9866 4240
rect 11282 4092 11386 4240
rect 8653 4040 10975 4041
rect 8653 1720 8654 4040
rect 10974 1720 10975 4040
rect 8653 1719 10975 1720
rect 7784 1292 7888 1668
rect 5155 1240 7477 1241
rect 5155 -1080 5156 1240
rect 7476 -1080 7477 1240
rect 5155 -1081 7477 -1080
rect 4286 -1508 4390 -1132
rect 1657 -1560 3979 -1559
rect 1657 -3880 1658 -1560
rect 3978 -3880 3979 -1560
rect 1657 -3881 3979 -3880
rect 788 -4080 892 -3932
rect 2766 -4080 2870 -3881
rect 4286 -3932 4306 -1508
rect 4370 -3932 4390 -1508
rect 6264 -1559 6368 -1081
rect 7784 -1132 7804 1292
rect 7868 -1132 7888 1292
rect 9762 1241 9866 1719
rect 11282 1668 11302 4092
rect 11366 1668 11386 4092
rect 11282 1292 11386 1668
rect 8653 1240 10975 1241
rect 8653 -1080 8654 1240
rect 10974 -1080 10975 1240
rect 8653 -1081 10975 -1080
rect 7784 -1508 7888 -1132
rect 5155 -1560 7477 -1559
rect 5155 -3880 5156 -1560
rect 7476 -3880 7477 -1560
rect 5155 -3881 7477 -3880
rect 4286 -4080 4390 -3932
rect 6264 -4080 6368 -3881
rect 7784 -3932 7804 -1508
rect 7868 -3932 7888 -1508
rect 9762 -1559 9866 -1081
rect 11282 -1132 11302 1292
rect 11366 -1132 11386 1292
rect 11282 -1508 11386 -1132
rect 8653 -1560 10975 -1559
rect 8653 -3880 8654 -1560
rect 10974 -3880 10975 -1560
rect 8653 -3881 10975 -3880
rect 7784 -4080 7888 -3932
rect 9762 -4080 9866 -3881
rect 11282 -3932 11302 -1508
rect 11366 -3932 11386 -1508
rect 11282 -4080 11386 -3932
<< properties >>
string FIXED_BBOX 6144 1480 8624 3960
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 12 l 12 val 297.12 carea 2.00 cperi 0.19 class capacitor nx 6 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
